// Commented out to prevent synthesis issues
// `default_nettype none

module ChipInterface (  
    input  logic        CLOCK_100, // 100 MHz Clock
    output logic        i2s0_sck, i2s0_ws, 
    input  logic        i2s0_sd,
    output logic        i2s1_sck, i2s1_ws, 
    input  logic        i2s1_sd,
    output logic        uart0_tx,
    input  logic [15:0] SW,
    output logic [15:0] LD,
    input  logic [ 3:0] BTN,
    output logic [ 7:0] D0_SEG, D1_SEG,
    output logic [ 3:0] D0_AN, D1_AN
);

    import utils::*;

    logic [ 6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7;
    logic [31:0] BCD_LT, BCD_RT;

    SevenSegmentDisplay ssd (.BCD7(BCD_RT[15:12]),  
                             .BCD6(BCD_RT[11:8]),
                             .BCD5(BCD_RT[7:4]),
                             .BCD4(BCD_RT[3:0]),
                             .BCD3(BCD_LT[15:12]),
                             .BCD2(BCD_LT[11:8]),
                             .BCD1(BCD_LT[7:4]),
                             .BCD0(BCD_LT[3:0]),
                             .blank(8'b0),
                             .HEX7,
                             .HEX6,
                             .HEX5,
                             .HEX4,
                             .HEX3,
                             .HEX2,
                             .HEX1,
                             .HEX0);

    SSegDisplayDriver ssdd (.clk(CLOCK_100),
                            .reset(BTN[0]),
                            .HEX0,
                            .HEX1,
                            .HEX2,
                            .HEX3,
                            .HEX4,
                            .HEX5,
                            .HEX6,
                            .HEX7,
                            .dpoints(8'b0000_0000),
                            .D1_AN(D0_AN),
                            .D2_AN(D1_AN),
                            .D1_SEG(D0_SEG),
                            .D2_SEG(D1_SEG));

    logic [1:0][17:0] data;
    logic [1:0]       data_rdy;

    I2SInterface i2s0 (.clock(CLOCK_100),
                       .reset(BTN[0]),
                       .I2S_SCK(i2s0_sck),
                       .I2S_WS(i2s0_ws),
                       .I2S_SD(i2s0_sd),
                       .data(data[0]),
                       .d_rdy_l(data_rdy[0]),
                       .d_rdy_r());

    I2SInterface i2s1 (.clock(CLOCK_100),
                       .reset(BTN[0]),
                       .I2S_SCK(i2s1_sck),
                       .I2S_WS(i2s1_ws),
                       .I2S_SD(i2s1_sd),
                       .data(data[1]),
                       .d_rdy_l(data_rdy[1]),
                       .d_rdy_r());
    
    DisplaySamples #(.CALIB_VAL(13'd7296))
                rd0 (.clock(CLOCK_100),
                     .reset(BTN[0]),
                     .data(data[0]),
                     .data_rdy(data_rdy[0]),
                     .disp_val(BCD_LT));

    DisplaySamples #(.CALIB_VAL(13'd7040))
                rd1 (.clock(CLOCK_100),
                     .reset(BTN[0]),
                     .data(data[1]),
                     .data_rdy(data_rdy[1]),
                     .disp_val(BCD_RT));

    logic [1:0] noise_detected, start_calc;

    assign LD[ 7:0] = (noise_detected[0]) ? 8'b1111_1111 : 0;
    assign LD[15:8] = (noise_detected[1]) ? 8'b1111_1111 : 0;
    
    // Left mic
    // NOTE: buf 0 is our reference.
    // we're only running threshold detection on buf0, so we'll
    // cross-correlate it to buf1 and argmax on the shift to buf1 (k),
    // giving us k_hat, will be used as the index into the LUT.
    Buffer #(.THRESHOLD(13'd4_096), .CALIB_VAL(13'd7_296))
           buf0 (.clock(CLOCK_100),
                 .reset(BTN[0]),
                 .restart(BTN[1]),
                 .data_in(data[0]),
                 .data_rdy(data_rdy[0]),
                 .read_offset(addr0),
                 .finished_calc(tdoa_done),
                 .data_out(sample0),
                 .noise_detected(noise_detected[0]),
                 .start_calc(start_calc[0]));

    // Right mic
    Buffer #(.THRESHOLD(13'd4_096), .CALIB_VAL(13'd7_040))
           buf1 (.clock(CLOCK_100),
                 .reset(BTN[0]),
                 .restart(BTN[1]),
                 .data_in(data[1]),
                 .data_rdy(data_rdy[1]),
                 .read_offset(addr1),
                 .finished_calc(tdoa_done),
                 .data_out(sample1),
                 .noise_detected(noise_detected[1]),
                 .start_calc(start_calc[1]));

    TDOA tdoa (.clock(CLOCK_100),
               .reset(BTN[0]),
               .restart(BTN[1]),
               .ready(start_calc[0]),
               .din0(sample0),
               .din1(sample1),
               .addr0,
               .addr1,
               .done(tdoa_done), 
               .k_hat);

    blk_mem_gen_0 lut (.clka(CLOCK_100),
                       .addra(lut_idx),
                       .douta(angle));

    logic [8:0]  addr0, addr1;
    logic [17:0] sample0, sample1;
    logic [7:0]  k_hat, lut_idx;
    logic [7:0]  angle;
    logic        tdoa_done, tx_busy, angle_rdy;

    assign angle_rdy = tdoa_done & ~tx_busy;

    always_comb begin
        if (-k_hat > 8'd42) lut_idx = 0;
        else if (k_hat > 8'd42) lut_idx = 8'd84;
        else lut_idx = k_hat + 8'd42;
    end

    UARTInterface uart0 (.clock(CLOCK_100),
                         .reset(BTN[0]),
                         .data_rdy(angle_rdy),
                         .data(angle),
                         .UART_TX(uart0_tx),
                         .tx_busy);

endmodule : ChipInterface